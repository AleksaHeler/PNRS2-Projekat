interface device_if;
    
endinterface