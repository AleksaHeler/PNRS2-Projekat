//  Class: apb_sequencer
//
class apb_sequencer extends uvm_sequencer#(sequence_item);
    `uvm_component_utils(apb_sequencer);

    //  Group: Configuration Object(s)

    
    //  Group: Components


    //  Group: Variables


    //  Group: Functions

    //  Constructor: new
    function new(string name = "apb_sequencer", uvm_component parent);
        super.new(name, parent);
    endfunction: new

    
endclass: apb_sequencer
