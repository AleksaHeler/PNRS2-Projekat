package my_package;
   import uvm_pkg::*;
`include "uvm_macros.svh"

`include "coverage.sv"
`include "sequence_item.sv"
`include "sequencer.sv"
`include "sequence.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "environment.sv"
`include "basic_test.sv"
`include "wr_rd_test.sv"
`include "all_wr_rd_test.sv"
`include "deterministic_all_wr_rd_test.sv"

endpackage : my_package
  