package my_package;

`include "transaction.sv"

endpackage : my_package
  