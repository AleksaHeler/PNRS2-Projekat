class driver extends uvm_driver;

endclass